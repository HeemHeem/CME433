`ifndef PARAMETERS
`define T    3
`define LOW  5
`define MED  10
`define HIGH 15
`endif
