----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:33:16 10/08/2010 
-- Design Name: 
-- Module Name:    davio - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Parity_davio is
port (D   : in std_logic_vector(6 downto 0);
      F   : out std_logic);
end Parity_davio;

architecture Behavioral of Parity_davio is
signal f6_0 : std_logic;
signal f6_2 : std_logic;
signal f5_0 : std_logic;
signal f5_2 : std_logic;
begin
	f6_0 <=
	
	f6_2 <=

	f5_0 <=
			
	f5_2 <=
	
	F <=

end Behavioral;

